module pipeline_controller(
    input logic clk,
    input logic reset_n,
    input logic[4:0] rd,
    input logic[4:0] reg_1_addr,
    input logic[4:0] reg_2_addr,
    input logic new_rd,
    input logic reg_write,
    output logic forward
    
);

logic[4:0] past_rd;



endmodule 