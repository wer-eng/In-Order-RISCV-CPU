module hazard_unit(
    input logic jump,
    input logic branch,
    input logic[4:0] rd,
    output logic flush,
    output logic 

);


endmodule